-- Declaración de la entidad ---------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.componentes_pkg.all;

entity calculadora is
    port ();
end calculadora;

------ Arquitectura e Implementación de la Calculadora -----------
architecture arch of calculadora is

begin

end architecture;